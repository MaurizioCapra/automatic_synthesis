

module inv_beh( 
	input A,
	output Z);
	
	assign Z = !A;

endmodule
